module testbench();

reg q1, q2, q3, q4,q5, q6, q7, q8, q9, q10, q11, q12, q13, q14, q15, q16, q17, q18, q19, q20, q21, q22, q23, q24, q25, q26, q27, q28, q29, q30;
wire v1, v2, v3, v4, v5, v6, v7, v8;

tabla_1 U1(q1, q2, q3, v1);
tabla_2 U2(q4, q5, q6, v2);
tabla_3 U3(q7, q8, q9, q10, v3);
tabla_4 U4(q11, q12, q13, q14, v4);
tabla_5 U5(q15, q16, q17, q20, v5);
tabla_6 U6(q21, q22, q23, v6);
tabla_7 U7(q24, q25, q26, q27, v7);
tabla_8 U8(q28, q29, q30, v8);

initial begin
  #1
  $display("A B C | Y");
  $display("------|--");
  $monitor("%b %b %b | %b", q1, q2, q3, v1);
     q1 = 0; q2 = 0; q3 = 0;
  #1 q1 = 0; q2 = 0; q3 = 1;
  #1 q1 = 0; q2 = 1; q3 = 0;
  #1 q1 = 0; q2 = 1; q3 = 1;
  #1 q1 = 1; q2 = 0; q3 = 0;
  #1 q1 = 1; q2 = 0; q3 = 1;
  #1 q1 = 1; q2 = 1; q3 = 0;
  #1 q1 = 1; q2 = 1; q3 = 1;
end

initial begin
  #2
  $display("A B C | Y");
  $display("------|--");
  $monitor("%b %b %b | %b", q4, q5, q6, v2);
     q4 = 0; q5 = 0; q6 = 0;
  #1 q4 = 0; q5 = 0; q6 = 1;
  #1 q4 = 0; q5 = 1; q6 = 0;
  #1 q4 = 0; q5 = 1; q6 = 1;
  #1 q4 = 1; q5 = 0; q6 = 0;
  #1 q4 = 1; q5 = 0; q6 = 1;
  #1 q4 = 1; q5 = 1; q6 = 0;
  #1 q4 = 1; q5 = 1; q6 = 1;
end

initial begin
  #3
  $display("A B C D | Y");
  $display("--------|--");
  $monitor("%b %b %b %b | %b", q7, q8, q9, q10, v3);
     q7 = 0; q8 = 0; q9 = 0; q10 = 0;
  #1 q7 = 0; q8 = 0; q9 = 0; q10 = 1;
  #1 q7 = 0; q8 = 0; q9 = 1; q10 = 0;
  #1 q7 = 0; q8 = 0; q9 = 1; q10 = 1;
  #1 q7 = 0; q8 = 1; q9 = 0; q10 = 0;
  #1 q7 = 0; q8 = 1; q9 = 0; q10 = 1;
  #1 q7 = 0; q8 = 1; q9 = 1; q10 = 0;
  #1 q7 = 0; q8 = 1; q9 = 1; q10 = 1;
  #1 q7 = 1; q8 = 0; q9 = 0; q10 = 0;
  #1 q7 = 1; q8 = 0; q9 = 0; q10 = 1;
  #1 q7 = 1; q8 = 0; q9 = 1; q10 = 0;
  #1 q7 = 1; q8 = 0; q9 = 1; q10 = 1;
  #1 q7 = 1; q8 = 1; q9 = 0; q10 = 0;
  #1 q7 = 1; q8 = 1; q9 = 0; q10 = 1;
  #1 q7 = 1; q8 = 1; q9 = 1; q10 = 0;
  #1 q7 = 1; q8 = 1; q9 = 1; q10 = 1;

end

initial begin
  #4
  $display("A B C D | Y");
  $display("--------|--");
  $monitor("%b %b %b %b | %b", q11, q12, q13, q14, v4);
     q11 = 0; q12 = 0; q13 = 0; q14 = 0;
  #1 q11 = 0; q12 = 0; q13 = 0; q14 = 1;
  #1 q11 = 0; q12 = 0; q13 = 1; q14 = 0;
  #1 q11 = 0; q12 = 0; q13 = 1; q14 = 1;
  #1 q11 = 0; q12 = 1; q13 = 0; q14 = 0;
  #1 q11 = 0; q12 = 1; q13 = 0; q14 = 1;
  #1 q11 = 0; q12 = 1; q13 = 1; q14 = 0;
  #1 q11 = 0; q12 = 1; q13 = 1; q14 = 1;
  #1 q11 = 1; q12 = 0; q13 = 0; q14 = 0;
  #1 q11 = 1; q12 = 0; q13 = 0; q14 = 1;
  #1 q11 = 1; q12 = 0; q13 = 1; q14 = 0;
  #1 q11 = 1; q12 = 0; q13 = 1; q14 = 1;
  #1 q11 = 1; q12 = 1; q13 = 0; q14 = 0;
  #1 q11 = 1; q12 = 1; q13 = 0; q14 = 1;
  #1 q11 = 1; q12 = 1; q13 = 1; q14 = 0;
  #1 q11 = 1; q12 = 1; q13 = 1; q14 = 1;

end
///// ejercicio 2
initial begin
  #1
  $display("A B C D | Y");
  $display("--------|--");
  $monitor("%b %b %b %b | %b", q15, q16, q17, q20, v5);
     q15 = 0; q16 = 0; q17 = 0; q20 = 0;
  #1 q15 = 0; q16 = 0; q17 = 0; q20 = 1;
  #1 q15 = 0; q16 = 0; q17 = 1; q20 = 0;
  #1 q15 = 0; q16 = 0; q17 = 1; q20 = 1;
  #1 q15 = 0; q16 = 1; q17 = 0; q20 = 0;
  #1 q15 = 0; q16 = 1; q17 = 0; q20 = 1;
  #1 q15 = 0; q16 = 1; q17 = 1; q20 = 0;
  #1 q15 = 0; q16 = 1; q17 = 1; q20 = 1;
  #1 q15 = 1; q16 = 0; q17 = 0; q20 = 0;
  #1 q15 = 1; q16 = 0; q17 = 0; q20 = 1;
  #1 q15 = 1; q16 = 0; q17 = 1; q20 = 0;
  #1 q15 = 1; q16 = 0; q17 = 1; q20 = 1;
  #1 q15 = 1; q16 = 1; q17 = 0; q20 = 0;
  #1 q15 = 1; q16 = 1; q17 = 0; q20 = 1;
  #1 q15 = 1; q16 = 1; q17 = 1; q20 = 0;
  #1 q15 = 1; q16 = 1; q17 = 1; q20 = 1;

end

initial begin
  #2
  $display("A B C | Y");
  $display("------|--");
  $monitor("%b %b %b | %b", q21, q22, q23, v6);
     q21 = 0; q22 = 0; q23 = 0;
  #1 q21 = 0; q22 = 0; q23 = 1;
  #1 q21 = 0; q22 = 1; q23 = 0;
  #1 q21 = 0; q22 = 1; q23 = 1;
  #1 q21 = 1; q22 = 0; q23 = 0;
  #1 q21 = 1; q22 = 0; q23 = 1;
  #1 q21 = 1; q22 = 1; q23 = 0;
  #1 q21 = 1; q22 = 1; q23 = 1;
end

initial begin
  #3
  $display("A B C D | Y");
  $display("--------|--");
  $monitor("%b %b %b %b | %b", q24, q25, q26, q27, v7);
     q24 = 0; q25 = 0; q26 = 0; q27 = 0;
  #1 q24 = 0; q25 = 0; q26 = 0; q27 = 1;
  #1 q24 = 0; q25 = 0; q26 = 1; q27 = 0;
  #1 q24 = 0; q25 = 0; q26 = 1; q27 = 1;
  #1 q24 = 0; q25 = 1; q26 = 0; q27 = 0;
  #1 q24 = 0; q25 = 1; q26 = 0; q27 = 1;
  #1 q24 = 0; q25 = 1; q26 = 1; q27 = 0;
  #1 q24 = 0; q25 = 1; q26 = 1; q27 = 1;
  #1 q24 = 1; q25 = 0; q26 = 0; q27 = 0;
  #1 q24 = 1; q25 = 0; q26 = 0; q27 = 1;
  #1 q24 = 1; q25 = 0; q26 = 1; q27 = 0;
  #1 q24 = 1; q25 = 0; q26 = 1; q27 = 1;
  #1 q24 = 1; q25 = 1; q26 = 0; q27 = 0;
  #1 q24 = 1; q25 = 1; q26 = 0; q27 = 1;
  #1 q24 = 1; q25 = 1; q26 = 1; q27 = 0;
  #1 q24 = 1; q25 = 1; q26 = 1; q27 = 1;

end

initial begin
  #4
  $display("A B C | Y");
  $display("------|--");
  $monitor("%b %b %b | %b", q28, q29, q30, v8);
     q28 = 0; q29 = 0; q30 = 0;
  #1 q28 = 0; q29 = 0; q30 = 1;
  #1 q28 = 0; q29 = 1; q30 = 0;
  #1 q28 = 0; q29 = 1; q30 = 1;
  #1 q28 = 1; q29 = 0; q30 = 0;
  #1 q28 = 1; q29 = 0; q30 = 1;
  #1 q28 = 1; q29 = 1; q30 = 0;
  #1 q28 = 1; q29 = 1; q30 = 1;
end

initial
  #1 $finish;

initial begin
  $dumpfile("1.1_tb.vcd");
  $dumpvars(0, testbench);
end

endmodule




